module midi_freq_lut (
    input [6:0] note,
    output reg [23:0] frequency_x1000
);
    always @(*) begin
        case (note)
            7'd0: frequency_x1000 = 24'd8176;
            7'd1: frequency_x1000 = 24'd8662;
            7'd2: frequency_x1000 = 24'd9177;
            7'd3: frequency_x1000 = 24'd9723;
            7'd4: frequency_x1000 = 24'd10301;
            7'd5: frequency_x1000 = 24'd10913;
            7'd6: frequency_x1000 = 24'd11562;
            7'd7: frequency_x1000 = 24'd12250;
            7'd8: frequency_x1000 = 24'd12978;
            7'd9: frequency_x1000 = 24'd13750;
            7'd10: frequency_x1000 = 24'd14568;
            7'd11: frequency_x1000 = 24'd15434;
            7'd12: frequency_x1000 = 24'd16352;
            7'd13: frequency_x1000 = 24'd17324;
            7'd14: frequency_x1000 = 24'd18354;
            7'd15: frequency_x1000 = 24'd19445;
            7'd16: frequency_x1000 = 24'd20602;
            7'd17: frequency_x1000 = 24'd21827;
            7'd18: frequency_x1000 = 24'd23125;
            7'd19: frequency_x1000 = 24'd24500;
            7'd20: frequency_x1000 = 24'd25957;
            7'd21: frequency_x1000 = 24'd27500;
            7'd22: frequency_x1000 = 24'd29135;
            7'd23: frequency_x1000 = 24'd30868;
            7'd24: frequency_x1000 = 24'd32703;
            7'd25: frequency_x1000 = 24'd34648;
            7'd26: frequency_x1000 = 24'd36708;
            7'd27: frequency_x1000 = 24'd38891;
            7'd28: frequency_x1000 = 24'd41203;
            7'd29: frequency_x1000 = 24'd43654;
            7'd30: frequency_x1000 = 24'd46249;
            7'd31: frequency_x1000 = 24'd48999;
            7'd32: frequency_x1000 = 24'd51913;
            7'd33: frequency_x1000 = 24'd55000;
            7'd34: frequency_x1000 = 24'd58270;
            7'd35: frequency_x1000 = 24'd61735;
            7'd36: frequency_x1000 = 24'd65406;
            7'd37: frequency_x1000 = 24'd69296;
            7'd38: frequency_x1000 = 24'd73416;
            7'd39: frequency_x1000 = 24'd77782;
            7'd40: frequency_x1000 = 24'd82407;
            7'd41: frequency_x1000 = 24'd87307;
            7'd42: frequency_x1000 = 24'd92499;
            7'd43: frequency_x1000 = 24'd97999;
            7'd44: frequency_x1000 = 24'd103826;
            7'd45: frequency_x1000 = 24'd110000;
            7'd46: frequency_x1000 = 24'd116541;
            7'd47: frequency_x1000 = 24'd123471;
            7'd48: frequency_x1000 = 24'd130813;
            7'd49: frequency_x1000 = 24'd138591;
            7'd50: frequency_x1000 = 24'd146832;
            7'd51: frequency_x1000 = 24'd155563;
            7'd52: frequency_x1000 = 24'd164814;
            7'd53: frequency_x1000 = 24'd174614;
            7'd54: frequency_x1000 = 24'd184997;
            7'd55: frequency_x1000 = 24'd195998;
            7'd56: frequency_x1000 = 24'd207652;
            7'd57: frequency_x1000 = 24'd220000;
            7'd58: frequency_x1000 = 24'd233082;
            7'd59: frequency_x1000 = 24'd246942;
            7'd60: frequency_x1000 = 24'd261626;
            7'd61: frequency_x1000 = 24'd277183;
            7'd62: frequency_x1000 = 24'd293665;
            7'd63: frequency_x1000 = 24'd311127;
            7'd64: frequency_x1000 = 24'd329628;
            7'd65: frequency_x1000 = 24'd349228;
            7'd66: frequency_x1000 = 24'd369994;
            7'd67: frequency_x1000 = 24'd391995;
            7'd68: frequency_x1000 = 24'd415305;
            7'd69: frequency_x1000 = 24'd440000;
            7'd70: frequency_x1000 = 24'd466164;
            7'd71: frequency_x1000 = 24'd493883;
            7'd72: frequency_x1000 = 24'd523251;
            7'd73: frequency_x1000 = 24'd554365;
            7'd74: frequency_x1000 = 24'd587330;
            7'd75: frequency_x1000 = 24'd622254;
            7'd76: frequency_x1000 = 24'd659255;
            7'd77: frequency_x1000 = 24'd698456;
            7'd78: frequency_x1000 = 24'd739989;
            7'd79: frequency_x1000 = 24'd783991;
            7'd80: frequency_x1000 = 24'd830609;
            7'd81: frequency_x1000 = 24'd880000;
            7'd82: frequency_x1000 = 24'd932328;
            7'd83: frequency_x1000 = 24'd987767;
            7'd84: frequency_x1000 = 24'd1046502;
            7'd85: frequency_x1000 = 24'd1108731;
            7'd86: frequency_x1000 = 24'd1174659;
            7'd87: frequency_x1000 = 24'd1244508;
            7'd88: frequency_x1000 = 24'd1318510;
            7'd89: frequency_x1000 = 24'd1396913;
            7'd90: frequency_x1000 = 24'd1479978;
            7'd91: frequency_x1000 = 24'd1567982;
            7'd92: frequency_x1000 = 24'd1661219;
            7'd93: frequency_x1000 = 24'd1760000;
            7'd94: frequency_x1000 = 24'd1864655;
            7'd95: frequency_x1000 = 24'd1975533;
            7'd96: frequency_x1000 = 24'd2093005;
            7'd97: frequency_x1000 = 24'd2217461;
            7'd98: frequency_x1000 = 24'd2349318;
            7'd99: frequency_x1000 = 24'd2489016;
            7'd100: frequency_x1000 = 24'd2637020;
            7'd101: frequency_x1000 = 24'd2793826;
            7'd102: frequency_x1000 = 24'd2959955;
            7'd103: frequency_x1000 = 24'd3135963;
            7'd104: frequency_x1000 = 24'd3322438;
            7'd105: frequency_x1000 = 24'd3520000;
            7'd106: frequency_x1000 = 24'd3729310;
            7'd107: frequency_x1000 = 24'd3951066;
            7'd108: frequency_x1000 = 24'd4186009;
            7'd109: frequency_x1000 = 24'd4434922;
            7'd110: frequency_x1000 = 24'd4698636;
            7'd111: frequency_x1000 = 24'd4978032;
            7'd112: frequency_x1000 = 24'd5274041;
            7'd113: frequency_x1000 = 24'd5587652;
            7'd114: frequency_x1000 = 24'd5919911;
            7'd115: frequency_x1000 = 24'd6271927;
            7'd116: frequency_x1000 = 24'd6644875;
            7'd117: frequency_x1000 = 24'd7040000;
            7'd118: frequency_x1000 = 24'd7458620;
            7'd119: frequency_x1000 = 24'd7902133;
            7'd120: frequency_x1000 = 24'd8372018;
            7'd121: frequency_x1000 = 24'd8869844;
            7'd122: frequency_x1000 = 24'd9397273;
            7'd123: frequency_x1000 = 24'd9956063;
            7'd124: frequency_x1000 = 24'd10548082;
            7'd125: frequency_x1000 = 24'd11175303;
            7'd126: frequency_x1000 = 24'd11839822;
            7'd127: frequency_x1000 = 24'd12543854;
            default: frequency_x1000 = 24'd0;
        endcase
    end
endmodule
